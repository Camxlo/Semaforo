library verilog;
use verilog.vl_types.all;
entity Mod_Nocturno_vlg_vec_tst is
end Mod_Nocturno_vlg_vec_tst;
